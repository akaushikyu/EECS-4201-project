/*
 * Module: pd1
 *
 * Description: Top level module that will contain sub-module instantiations. 
 *
 * Inputs:
 * 1) clk
 * 2) reset signal
 */

module pd1 #(
    parameter int AWIDTH = 32,
    parameter int DWIDTH = 32)(
    input logic clk,
    input logic reset
);

 /*
  * Instantiate other submodules and 
  * probes. To be filled by student...
  *
  */



endmodule : pd1
