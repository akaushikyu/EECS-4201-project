mo@MoPC-Arch.73304:1768277015