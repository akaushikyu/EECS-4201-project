// ----  Probes  ----
`define PROBE_ASSIGN_XOR_OP1 assign_xor_op1
`define PROBE_ASSIGN_XOR_OP2 assign_xor_op2
`define PROBE_ASSIGN_XOR_RES assign_xor_res

// Define other probes as required....
`define ALU_OP1
`define ALU_OP2
`define ALU_RES
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd0 
// ----  Top module  ----
