/*
 *
 Module: three_stage_pipeline
 *
 * A 3-stage pipeline (TSP) where the first stage performs an addition of two
 * operands (op1_i, op2_i) and registers the output, and the second stage computes
 * the difference between the output from the first stage and op1_i and registers the
 * output. This means that the output (res_o) must be available two cycles after the
 * corresponding inputs have been observed on the rising clock edge
 *
 * Visually, the circuit should look like this:
 *               <---         Stage 1           --->
 *                                                        <---         Stage 2           --->
 *                                                                                               <--    Stage 3    -->
 *                                    |------------------>|                    |
 * -- op1_i -->|                    | --> |         |     |                    |-->|         |   |                    |
 *             | pipeline registers |     | ALU add | --> | pipeline registers |   | ALU sub |-->| pipeline register  | -- res_o -->
 * -- op2_i -->|                    | --> |         |     |                    |-->|         |   |                    |
 *
 * Inputs:
 * 1) 1-bit clock signal
 * 2) 1-bit wide synchronous reset
 * 3) DWIDTH-wide input op1_i
 * 4) DWIDTH-wide input op2_i
 *
 * Outputs:
 * 1) DWIDTH-wide result res_o
 */



import alu::*;
import reg_rst::*;

module three_stage_pipeline #(
			                  parameter int DWIDTH = 8)(
			                                            input logic               clk,
			                                            input logic               rst,
			                                            input logic [DWIDTH-1:0]  op1_i,
			                                            input logic [DWIDTH-1:0]  op2_i,
			                                            output logic [DWIDTH-1:0] res_o
			                                            );

  /*
   * Process definitions to be filled by
   * student below...
   * [HINT] Instantiate the alu and reg_rst modules
   * and set up the necessary connections
   *
   */
  int dwx2 = DWIDTH*2; 
  wire [DWIDTH*2-1:0] inS1;   wire [DWIDTH*2-1:0]inS1;

  wire [DWIDTH*2-1:0]inS1;
  wire [DWIDTH*2-1:0] inAluAdd;
  wire [DWIDTH*2-1:0] inAluSub;
  
  assign inS1[DWIDTH-1:0] = op1_i; 
  assign inS1[DWIDTH*2-1:DWIDTH] = op2_i;
  
  wire [DWIDTH*2-1:0]inS2;
  wire [DWIDTH-1:0]  outAluAdd;
  wire [DWIDTH-1:0]  outAluSub;
  
  assign inS2[DWIDTH*2-1:0] = op1_i + (outAluAdd << (DWIDTH-1));
  
  wire [DWIDTH-1:0]inS3;
  
  reg_rst #(.dwx2) s1(.clk(clk),.rst(rst),.in_i(inS1),.out_i(inAluAdd));
  reg_rst #(.dwx2) s2(.clk(clk),.rst(rst),.in_i(inS1[DWIDTH-1:0]+(outAluAdd<<(DWIDTH-1))),.out_i(inS2)); 
  reg_rst #(.dwx2) s3(.clk(clk),.rst(rst),.in_i(outAluSub),.out_i(1'd0 + (inS3<<(DWIDTH-1))));	  
  alu #(.DWIDTH) adder(.clk(clk),.rst(rst),.op1_i(inAluAdd[DWIDTH*2-1:DWIDTH]),.op2_i(inAluAdd[DWIDTH-1:0]),.res_o(outAluAdd));
  alu #(.DWIDTH) subber(.clk(clk),.rst(rst),.op1_i(inAluSub[DWIDTH*2-1:DWIDTH]),.op2_i(inAluSub[DWIDTH-1:0]),.res_o(outAluSub));

  assign res_o = inS3[DWIDTH*2-1:DWIDTH];
  
  
  
  
endmodule: three_stage_pipeline
