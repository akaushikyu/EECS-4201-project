// ----  Probes  ----
//`define PROBE_F_PC // ??
//`define PROBE_F_INSN // ??

//`define PROBE_D_PC // ??
//`define PROBE_D_OPCODE // ??
//`define PROBE_D_RD // ??
//`define PROBE_D_FUNCT3 // ??
//`define PROBE_D_RS1 // ??
//`define PROBE_D_RS2 // ??
//`define PROBE_D_FUNCT7 // ??
//`define PROBE_D_IMM // ??
//`define PROBE_D_SHAMT // ??

//`define R_WRITE_ENABLE      // ??
//`define R_WRITE_DESTINATION // ??
//`define R_WRITE_DATA        // ??
//`define R_READ_RS1          // ??
//`define R_READ_RS2          // ??
//`define R_READ_RS1_DATA     // ??
//`define R_READ_RS2_DATA     // ??

//`define E_PC                // ??
//`define E_ALU_RES           // ??
//`define E_BR_TAKEN          // ??
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd3
// ----  Top module  ----
