/*
 * Module: igen
 *
 * Description: Immediate value generator
 * 
 * Inputs:
 * 1) opcode opcode_i
 * Outputs:
 * 2) 32-bit immediate value imm_o
 */

module igen (
    input logic [6:0] opcode_i,
    output logic [31:0] imm_o
);
    /*
     * Process definitions to be filled by 
     * student below...
     */

endmodule : igen
