// ----  Probes  ----
`define PROBE_ADDR      // ??
`define PROBE_DATA_IN   // ??
`define PROBE_DATA_OUT  // ??
`define PROBE_READ_EN   // ??
`define PROBE_WRITE_EN  // ??
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1 
// ----  Top module  ----
